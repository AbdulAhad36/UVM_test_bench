interface my_interface();

//inputs and  outputs

endinterface
